class yapp_tx_agent extends uvm_agent;
    `uvm_component_utils_begin(yapp_tx_agent)
    `uvm_field_enum(uvm_active_passive_enum, is_active, UVM_ALL_ON)
    `uvm_component_utils_end
    function new(string name, uvm_component parent);
        super.new(name, parent);
    endfunction

    yapp_tx_driver driver;
    yapp_tx_monitor monitor;
    yapp_tx_sequencer sequencer;

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        monitor = new("monitor", this);
        if(is_active == UVM_ACTIVE) begin
            sequencer = new("sequencer", this);
            driver = new("driver", this);
        end
    endfunction

    function void connect_phase(uvm_phase phase);
        if(is_active == UVM_ACTIVE) begin
            driver.seq_item_port.connect(sequencer.seq_item_export);
        end
    endfunction

    function void start_of_simulation_phase(uvm_phase phase);
        `uvm_info(get_type_name(),"Running Simulation...", UVM_HIGH);
    endfunction

endclass